module sound

pub struct Sound {
mut:
	path string
	volume f32
	x f32
	z f32
}