module sound

pub struct SoundEngine {
	
}