module components

pub struct Location {
mut:
	x f32
	y f32
}